`timescale 1ns / 1ps
`define period 10
////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:57:40 08/12/2017
// Design Name:   Ray_AABB_32bit
// Module Name:   C:/Users/George/Dropbox/Imperial_College_London/Thesis/RTL/flopoco/Ray_AABB_11_52_pipelined_correctR/tb11_52.v
// Project Name:  Ray_AABB_11_52_pipelined_correctR
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Ray_AABB_32bit
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb11_52;

	// Inputs
	reg clk;
	reg rst;
	reg [65:0] x0UP;
	reg [65:0] x0LOW;
	reg [65:0] y0UP;
	reg [65:0] y0LOW;
	reg [65:0] z0UP;
	reg [65:0] z0LOW;
	reg [65:0] x1LOW;
	reg [65:0] y1LOW;
	reg [65:0] z1LOW;
	reg [65:0] x2UP;
	reg [65:0] y2UP;
	reg [65:0] z2UP;
	reg x;
	reg y;
	reg z;
	reg [65:0] divxUP;
	reg [65:0] divxLOW;
	reg [65:0] divyUP;
	reg [65:0] divyLOW;
	reg [65:0] divzUP;
	reg [65:0] divzLOW;

	// Outputs
	wire hit_miss;

	// Instantiate the Unit Under Test (UUT)
	Ray_AABB_11_52 uut (
		.clk(clk), 
		.rst(rst), 
		.x0UP(x0UP), 
		.x0LOW(x0LOW), 
		.y0UP(y0UP), 
		.y0LOW(y0LOW), 
		.z0UP(z0UP), 
		.z0LOW(z0LOW), 
		.x1LOW(x1LOW), 
		.y1LOW(y1LOW), 
		.z1LOW(z1LOW), 
		.x2UP(x2UP), 
		.y2UP(y2UP), 
		.z2UP(z2UP), 
		.x(x), 
		.y(y), 
		.z(z), 
		.divxUP(divxUP), 
		.divxLOW(divxLOW), 
		.divyUP(divyUP), 
		.divyLOW(divyLOW), 
		.divzUP(divzUP), 
		.divzLOW(divzLOW), 
		.hit_miss(hit_miss)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 1;
	
		x0UP = 66'b010011111111100110101101111111000110101001001001010010011111011000;
      x0LOW =66'b010011111111100110101101111111000110101001001001010010011111011000;
		y0UP = 66'b010011111111010011100010100100101001011011110000111100101100011011;
		y0LOW =66'b010011111111010011100010100100101001011011110000111100101100011011;
		z0UP = 66'b010011111111000100001001111010110110000011100001100101110011010001;
		z0LOW =66'b010011111111000100001001111010110110000011100001100101110011010001;
		x1LOW =66'b010011111110111011100001101001110110010011011110010100010000001111;

		y1LOW =66'b010011111110110011101010011001000011011101100010000101101111011010;

		z1LOW =66'b011011111111011101011111110110100000101010100010111100010011000101;

		x2UP = 66'b010011111111011101011110010000100000101001100110100010110100111101;

		y2UP = 66'b010011111111001011010010101000100110111100000000001111011110100010;

		z2UP = 66'b011011111110101101010101111001000101100001011001101100110100111111;

		x = 0;
		y = 0;
		z = 0;
		divxUP =66'b011011111111111000011001010111111000001001000110100101101011110101;
		divxLOW=66'b011011111111111000011001010111111000001001000110100101101011110101;
		divyUP =66'b011100000000001111110011000100110011011111101011001010001101100010;
		divyLOW=66'b011100000000001111110011000100110011011111101011001010001101100010;
		divzUP =66'b011011111111110101011010101001001100000000111110010010010001000100;
		divzLOW=66'b011011111111110101011010101001001100000000111110010010010001000100;

		#2;
		//#0.6916;
		rst = 0;
		
		#8
		//#2.7664;
		x0UP = 66'b011011111111100110111000011011111100000010000010001110111010111100; //hit2
		x0LOW = 66'b011011111111100110111000011011111100000010000010001110111010111100;
		y0UP = 66'b010011111110100110001111101000010011001011000000000110111011100110;
		y0LOW = 66'b010011111110100110001111101000010011001011000000000110111011100110;
		z0UP = 66'b010011111111011011101000011000110110000011111000011010000101110000;
		z0LOW = 66'b010011111111011011101000011000110110000011111000011010000101110000;
		x1LOW = 66'b011011111111101000110100011110011110011110100010100100010000111100;
		y1LOW = 66'b010011111110111010100111100110000011111110100111010111111101010111;
		z1LOW = 66'b010011111111100110111000111110100110110100011001000010000000111011;
		x2UP = 66'b011011111110101001000100100011111001000110000010111101001011110010;
		y2UP = 66'b010011111111100110110011001100101010110011111011011101100010110110;
		z2UP = 66'b010011111111100111100110100110110000100111011100001000011101010010;
		x = 0;
		y = 0;
		z = 0;
		divxUP = 66'b010100000000000010100101100001000001000010011011010110001011011010;
		divxLOW = 66'b010100000000000010100101100001000001000010011011010110001011011010;
		divyUP = 66'b010011111111110001011000110111010001011110011101101010110111011100;
		divyLOW = 66'b010011111111110001011000110111010001011110011101101010110111011100;
		divzUP = 66'b010011111111110011000111111110101011101100011100101000010010000010;
		divzLOW = 66'b010011111111110011000111111110101011101100011100101000010010000010;
		
		end
      always #(`period/2) clk = ~clk;
endmodule