`timescale 1ns / 1ps
`define period 10
////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:16:43 08/14/2017
// Design Name:   Ray_AABB_11_23
// Module Name:   C:/Users/George/Dropbox/Imperial_College_London/Thesis/RTL/flopoco/Ray_AABB_11_23_correctR/tb.v
// Project Name:  Ray_AABB_11_23_correctR
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Ray_AABB_11_23
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	reg clk;
	reg rst;
	reg [36:0] x0;
	reg [36:0] y0;
	reg [36:0] z0;
	reg [36:0] x1;
	reg [36:0] y1;
	reg [36:0] z1;
	reg [36:0] x2;
	reg [36:0] y2;
	reg [36:0] z2;
	reg [36:0] divx;
	reg [36:0] divy;
	reg [36:0] divz;
	reg x;
	reg y;
	reg z;
	// Outputs
	wire hit_miss;

	// Instantiate the Unit Under Test (UUT)
	Ray_AABB_11_23 uut (
		.clk(clk), 
		.rst(rst), 
		.x0(x0),  
		.y0(y0), 
		.z0(z0), 
		.x1(x1), 
		.y1(y1), 
		.z1(z1), 
		.x2(x2), 
		.y2(y2), 
		.z2(z2),  
		.divx(divx), 
		.divy(divy), 
		.divz(divz), 
		.x(x), 
		.y(y), 
		.z(z),
		.hit_miss(hit_miss)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 1;
		
      x0 = 37'b0100111111111001101011011111110001101;//hit1
		y0 = 37'b0100111111110100111000101001001010010;
		z0 = 37'b0100111111110001000010011110101101100;

		x1 = 37'b0100111111101110111000011010011101100;
		y1 = 37'b0100111111101100111010100110010000110;
		z1 = 37'b0110111111110111010111111101101000001;

		x2 = 37'b0100111111110111010111100100001000001;
		y2 = 37'b0100111111110010110100101010001001101;
		z2 = 37'b0110111111101011010101011110010001011;

		x = 0;
		y = 0;
		z = 0;
		divx = 37'b0110111111111110000110010101111110000;
		divy = 37'b0111000000000011111100110001001100110;
		divz = 37'b0110111111111101010110101010010011000;
		
		#2;
		//#0.6916;
		rst = 0;
		
		#8;
		//#2.7664;
		x0 = 37'b0110111111111010010001001110011000101; //hit3
		y0 = 37'b0100111111111000100001101010110110010;
		z0 = 37'b0110111111111001000111111011010110101;
		x1 = 37'b0110111111111001001010000001110111100;
		y1 = 37'b0110111111110110001111011010000010110;
		z1 = 37'b0110111111111011000111101100100010101;
		x2 = 37'b0100111111110001010101000010011111001;
		y2 = 37'b0100111111110000001110011000111100110;
		z2 = 37'b0110111111110010001100000011111001011;

		x = 0;
		y = 0;
		z = 0;       
		divx = 37'b0101000000000010111000110011101010101;
		divy = 37'b0110111111111101100000101000111111000;
		divz = 37'b0111000000000111001000101000011110111;
		
		#10;
		x0 = 37'b0100111111111001101011011111110001101; //hit-->miss
		y0 = 37'b0100111111110100111000101001001010010;
		z0 = 37'b0100111111110001000010011110101101100;
		x1 = 37'b0100111111101110111000011010011101100;
		y1 = 37'b0100111111101100111010100110010000110;
		z1 = 37'b0110111111110111010111111101101000001;
		x2 = 37'b0100111111110111010111100100001000001;
		y2 = 37'b0100111111110010110100101010001001101;
		z2 = 37'b0110111111101011010101011110010001011;
		x = 1;
		y = 0;
		z = 0;
		divx = 37'b0110111111111110000110010101111110000;
		divy = 37'b0111000000000011111100110001001100110;
		divz = 37'b0110111111111101010110101010010011000;

		#10;
		x0 = 37'b0110111111111001101110000110111111000; //hit2
		y0 = 37'b0100111111101001100011111010000100110;
		z0 = 37'b0100111111110110111010000110001101100;
		x1 = 37'b0110111111111010001101000111100111100;
		y1 = 37'b0100111111101110101001111001100000111;
		z1 = 37'b0100111111111001101110001111101001101;
		x2 = 37'b0110111111101010010001001000111110010;
		y2 = 37'b0100111111111001101100110011001010101;
		z2 = 37'b0100111111111001111001101001101100001;
		x = 0;
		y = 0;
		z = 0;
		divx = 37'b0101000000000000101001011000010000010;
		divy = 37'b0100111111111100010110001101110100010;
		divz = 37'b0100111111111100110001111111101010111;
		
		
		#10;
	//	#3.458;
      x0 = 37'b0110111111010111111001101110011100000; //miss
		y0 = 37'b0100111110110011101110000001101001000;
		z0 = 37'b0110111111011110100000010110000011000;
		x1 = 37'b0110111111011100010111110000000010000;
		y1 = 37'b0110111110110011111001110010100101000;
		z1 = 37'b0110111101111011101011111010110000000;
		x2=  37'b0110111111000000111100010100010111000;
		y2 = 37'b0100111111000001011010011011011001000;
		z2 = 37'b0100111111010110011111111110010010000;
		x = 0;
		y = 0;
		z = 0;
		divx = 37'b0100111111100001000110110010011010000;
		divy = 37'b0111000000001101010100110000010000000;
		divz = 37'b0110111111111011000010101001110010000;
	
		end
	
	always #(`period/2) clk = ~clk;
      
endmodule

